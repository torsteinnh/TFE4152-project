* This file contains the parameters and standard components for all analog circuits in the project.

* Include models

* Test parameters
.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]


* Derived and fixed test parameters
.param VDD = 1.8 ! Supply voltage
.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param READ_TIME = {CLK_PERIOD}
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param NRE_R2_DLY = {CLK_PERIOD + NRE_R1_DLY + READ_TIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {CLK_PERIOD + NRE_R2_DLY + READ_TIME} ! Delay for ERASE signal
.param PERIOD = {ERASE_DLY + EXPOSURETIME} ! Period for testbench sources


* Permanent test sources
VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF READ_TIME PERIOD)
VNRE_R2 NRE_R2 0 dc 0  pulse(VDD 0 NRE_R2_DLY TRF TRF READ_TIME PERIOD)


* Parameters for photo cell, L [0.36 , 1.08]u W [1.08 , 5.04]u
.param M1W = 1.08u
.param M1L = 1.08u
.param M2W = 1.08u
.param M2L = 1.08u
.param M3W = 3u
.param M3L = 0.67u
.param M4W = 1.08u
.param M4L = 1.08u
.param MCW = 1u
.param MCL = 1u

.param CSval = 2p
.param CCval = 3p
